//-----------------------------------------------------
// File Name   : alucodes.sv
// Function    : pMIPS ALU function code definitions 
// Author:   tjk
// Last rev. 23 Oct 12 
//-----------------------------------------------------
// 
`define RA   3'b000
`define RB   3'b001
`define RADD  3'b010
`define RSUB  3'b011  
`define RAND  3'b100
`define ROR   3'b101 
// `define RXOR  3'b110  
`define RNOP  3'b110  
// `define RNOR  3'b111
`define RMUL  3'b111